module name(a,b,c,x,y);

  output x,y;
  input a,b,c;

  //the body

endmodule;
